** Generated for: hspiceD
** Generated on: Nov 13 23:10:06 2022
** Design library name: mylib2
** Design cell name: myFATestbench
** Design view name: schematic

.GLOBAL vdd!
.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/NMOS_VTL.inc"
.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/PMOS_VTL.inc"
.include "fulladder.pex.netlist.pex"

.subckt fulladder  A COUT CIN S B GND! VDD!
* 
* VDD!	VDD!
* GND!	GND!
* B	B
* S	S
* CIN	CIN
* COUT	COUT
* A	A
mXI17/MM0 N_NET058_XI17/MM0_d N_A_XI17/MM0_g N_GND!_XI17/MM0_s N_GND!_XI17/MM0_b
+ NMOS_VTL L=5e-08 W=9e-08 AD=1.17e-14 AS=1.35e-14 PD=4.4e-07 PS=4.8e-07
mXI16/MM0 N_NET06_XI16/MM0_d N_NET058_XI16/MM0_g N_GND!_XI17/MM0_s
+ N_GND!_XI17/MM0_b NMOS_VTL L=5e-08 W=9e-08 AD=1.08e-14 AS=1.35e-14 PD=4.2e-07
+ PS=4.8e-07
mXI15/MM0 N_COUT_XI15/MM0_d N_NET27_XI15/MM0_g N_GND!_XI15/MM0_s
+ N_GND!_XI17/MM0_b NMOS_VTL L=5e-08 W=9e-08 AD=1.44e-14 AS=1.44e-14 PD=5e-07
+ PS=5e-07
MM8 N_NET50_MM8_d N_NET27_MM8_g N_NET37_MM8_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=3.06e-14 AS=3.06e-14 PD=7e-07 PS=7e-07
MM5 N_NET37_MM8_s N_NET06_MM5_g N_GND!_MM5_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=3.06e-14 AS=3.06e-14 PD=7e-07 PS=7e-07
MM2 N_NET16_MM2_d N_NET06_MM2_g N_GND!_MM2_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=3.06e-14 PD=6e-07 PS=7e-07
MM6 N_NET37_MM6_d N_NET031_MM6_g N_GND!_MM5_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=3.06e-14 AS=3.06e-14 PD=7e-07 PS=7e-07
MM3 N_NET16_MM3_d N_NET031_MM3_g N_GND!_MM2_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=3.06e-14 AS=3.06e-14 PD=7e-07 PS=7e-07
MM7 N_NET37_MM6_d N_CIN_MM7_g N_GND!_MM7_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=3.06e-14 AS=5.31e-14 PD=7e-07 PS=1.06e-06
MM0 N_NET27_MM0_d N_CIN_MM0_g N_NET16_MM3_d N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=4.68e-14 AS=3.06e-14 PD=8.8e-07 PS=7e-07
MM12 NET64 N_NET06_MM12_g N_GND!_MM7_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=2.7e-07 AD=3.78e-14 AS=5.31e-14 PD=8.2e-07 PS=1.06e-06
MM1 N_NET27_MM0_d N_NET06_MM1_g NET26 N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=4.68e-14 AS=2.52e-14 PD=8.8e-07 PS=6.4e-07
MM11 NET49 N_NET031_MM11_g NET64 N_GND!_XI17/MM0_b NMOS_VTL L=5e-08 W=2.7e-07
+ AD=5.13e-14 AS=3.78e-14 PD=9.2e-07 PS=8.2e-07
MM4 NET26 N_NET031_MM4_g N_GND!_MM4_s N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07
MM10 N_NET50_MM10_d N_CIN_MM10_g NET49 N_GND!_XI17/MM0_b NMOS_VTL L=5e-08
+ W=2.7e-07 AD=5.4e-14 AS=5.13e-14 PD=9.4e-07 PS=9.2e-07
mXI14/MM0 N_S_XI14/MM0_d N_NET50_XI14/MM0_g N_GND!_XI14/MM0_s N_GND!_XI17/MM0_b
+ NMOS_VTL L=5e-08 W=9e-08 AD=1.44e-14 AS=1.44e-14 PD=5e-07 PS=5e-07
mXI18/MM0 N_NET031_XI18/MM0_d N_NET059_XI18/MM0_g N_GND!_XI18/MM0_s
+ N_GND!_XI17/MM0_b NMOS_VTL L=5e-08 W=9e-08 AD=1.17e-14 AS=1.44e-14 PD=4.4e-07
+ PS=5e-07
mXI19/MM0 N_NET059_XI19/MM0_d N_B_XI19/MM0_g N_GND!_XI18/MM0_s N_GND!_XI17/MM0_b
+ NMOS_VTL L=5e-08 W=9e-08 AD=9.9e-15 AS=1.44e-14 PD=4e-07 PS=5e-07
mXI17/MM1 N_NET058_XI17/MM1_d N_A_XI17/MM1_g N_VDD!_XI17/MM1_s N_VDD!_XI17/MM1_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
mXI16/MM1 N_NET06_XI16/MM1_d N_NET058_XI16/MM1_g N_VDD!_XI17/MM1_s
+ N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07
+ PS=6.6e-07
mXI15/MM1 N_COUT_XI15/MM1_d N_NET27_XI15/MM1_g N_VDD!_XI15/MM1_s
+ N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.88e-14
+ PD=6.8e-07 PS=6.8e-07
MM19 N_NET50_MM19_d N_NET27_MM19_g N_NET41_MM19_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=6.12e-14 AS=6.12e-14 PD=1.06e-06 PS=1.06e-06
MM15 N_NET20_MM15_d N_NET06_MM15_g N_VDD!_MM15_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=4.32e-14 AS=6.12e-14 PD=9.6e-07 PS=1.06e-06
MM20 N_NET41_MM19_s N_NET06_MM20_g N_VDD!_MM20_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=6.12e-14 AS=6.12e-14 PD=1.06e-06 PS=1.06e-06
MM18 N_NET20_MM18_d N_NET031_MM18_g N_VDD!_MM15_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=6.12e-14 AS=6.12e-14 PD=1.06e-06 PS=1.06e-06
MM21 N_NET41_MM21_d N_NET031_MM21_g N_VDD!_MM20_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=6.12e-14 AS=6.12e-14 PD=1.06e-06 PS=1.06e-06
MM14 N_NET27_MM14_d N_CIN_MM14_g N_NET20_MM18_d N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=9.36e-14 AS=6.12e-14 PD=1.24e-06 PS=1.06e-06
MM22 N_NET41_MM21_d N_CIN_MM22_g N_VDD!_MM22_s N_VDD!_XI17/MM1_b PMOS_VTL
+ L=5e-08 W=3.6e-07 AD=6.12e-14 AS=1.062e-13 PD=1.06e-06 PS=1.6e-06
MM17 N_NET27_MM14_d N_NET06_MM17_g NET062 N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=9.36e-14 AS=5.04e-14 PD=1.24e-06 PS=1e-06
MM23 NET065 N_NET06_MM23_g N_VDD!_MM22_s N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=1.062e-13 PD=1.36e-06 PS=1.6e-06
MM16 NET062 N_NET031_MM16_g N_VDD!_MM16_s N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=5.04e-14 AS=5.04e-14 PD=1e-06 PS=1e-06
MM24 NET066 N_NET031_MM24_g NET065 N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08 W=5.4e-07
+ AD=1.026e-13 AS=7.56e-14 PD=1.46e-06 PS=1.36e-06
MM25 N_NET50_MM25_d N_CIN_MM25_g NET066 N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=1.08e-13 AS=1.026e-13 PD=1.48e-06 PS=1.46e-06
mXI14/MM1 N_S_XI14/MM1_d N_NET50_XI14/MM1_g N_VDD!_XI14/MM1_s N_VDD!_XI17/MM1_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.88e-14 PD=6.8e-07 PS=6.8e-07
mXI18/MM1 N_NET031_XI18/MM1_d N_NET059_XI18/MM1_g N_VDD!_XI18/MM1_s
+ N_VDD!_XI17/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.34e-14 AS=2.88e-14
+ PD=6.2e-07 PS=6.8e-07
mXI19/MM1 N_NET059_XI19/MM1_d N_B_XI19/MM1_g N_VDD!_XI18/MM1_s N_VDD!_XI17/MM1_b
+ PMOS_VTL L=5e-08 W=1.8e-07 AD=1.98e-14 AS=2.88e-14 PD=5.8e-07 PS=6.8e-07
*
.include "fulladder.pex.netlist.FULLADDER.pxi"
*
.ends
*
*

** Library name: mylib2
** Cell name: fulladdertb
** View name: schematic
xfulladder a cout cin s b gnd! vdd! fulladder  
c1 s 0 100e-15
c0 cout 0 100e-15


