*half adder
.TEMP 25
.OPTIONS ACCURATE
.OPTIONS POST=2

* YOU SHOULD INCLUDE MODLE FILES
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/NMOS_VTL.inc"
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/PMOS_VTL.inc"


* YOU SHOULD INCLUDE YOUR NELIST
.INCLUDE halfadder.sp

* YOU SHOULD ADD LOAD CAPACITANCE

* YOU SHOULD GIVE INPUT PATTERNS FOR SIMULATING POWER 

.PARAM PERIOD = 20NS
.PARAM T0= 0.1NS
.PARAM T1= T0+PERIOD
.PARAM T2= T1+0.1NS
.PARAM STEP= 1PS

*REPLACE "10NS" IN THE NEXT LINE WITH THE MEASURED WORST CASE DELAY OF YOUR OWN DESIGN
.PARAM DELAY_MAX= 0.7359NS

VDD   VDD! 0 0.7
VGND  GND! 0 0
.TRAN STEP T2

.MEASURE TOT_POWER AVG POWER FROM T0 TO T1

* THE POWER AT MAX FREQUENCY CAN BE CALCULATED BY DIVIDING THE SWITCHING ENERGY BY THE SWITCHING TIME
* YOU ONLY NEED TO REPORT THE POWER_AT_MAX VALUE. YOU DON'T NEED TO REPORT THE TOT_POWER VALUE
.MEASURE POWER_AT_MAX PARAM='TOT_POWER*PERIOD/DELAY_MAX'

.END








