*half adder
.TEMP 25
.OPTIONS ACCURATE
.OPTIONS POST=2

* YOU SHOULD INCLUDE MODLE FILES
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/NMOS_VTL.inc"
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/PMOS_VTL.inc"

* YOU SHOULD INCLUDE YOUR NELIST
.INCLUDE halfadder.sp

* YOU SHOULD ADD LOAD CAPACITANCE

* YOU SHOULD GIVE INPUT PATTERNS FOR TEST CASES
*Vin1 A gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 10n)
*Vin2 B gnd PULSE (0v 0.7v 9.9n 0.1n 0.1n 9.9n 20n)

* YOU SHOULD GIVE PROPER INPUT PATTERNS FOR MAXIMUM DELAY

.PARAM PERIOD = 20NS
.PARAM T0= 0.1NS
.PARAM T1= T0+PERIOD
.PARAM T2= T1+0.1NS
.PARAM STEP= 1PS

VDD   VDD! 0 0.7
VGND  GND! 0 0

.TRAN STEP T2

* YOU SHOULD MAKE SURE THAT YOU ARE MEASURING THE CORRECT SIGNAL FOR MAXIMUM DELAY. BELOW IS JUST AN EXAMPLE.
*.MEASURE TRAN DELAY_COUT1 TRIG V(a) VAL=0.35 RISE=1 TARG V(COUT) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_COUT2 TRIG V(a) VAL=0.35 RISE=1 TARG V(COUT) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_COUT3 TRIG V(a) VAL=0.35 FALL=1 TARG V(COUT) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_COUT4 TRIG V(a) VAL=0.35 FALL=1 TARG V(COUT) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_COUT5 TRIG V(b) VAL=0.35 RISE=1 TARG V(COUT) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_COUT6 TRIG V(b) VAL=0.35 RISE=1 TARG V(COUT) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_COUT7 TRIG V(b) VAL=0.35 FALL=1 TARG V(COUT) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_COUT8 TRIG V(b) VAL=0.35 FALL=1 TARG V(COUT) VAL= 0.35 FALL=1

*.MEASURE TRAN DELAY_S1 TRIG V(a) VAL=0.35 RISE=1 TARG V(S) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_S2 TRIG V(a) VAL=0.35 RISE=1 TARG V(S) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_S3 TRIG V(a) VAL=0.35 FALL=1 TARG V(S) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_S4 TRIG V(a) VAL=0.35 FALL=1 TARG V(S) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_S5 TRIG V(b) VAL=0.35 RISE=1 TARG V(S) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_S6 TRIG V(b) VAL=0.35 RISE=1 TARG V(S) VAL= 0.35 FALL=1
*.MEASURE TRAN DELAY_S7 TRIG V(b) VAL=0.35 FALL=1 TARG V(S) VAL= 0.35 RISE=1
*.MEASURE TRAN DELAY_S8 TRIG V(b) VAL=0.35 FALL=1 TARG V(S) VAL= 0.35 FALL=1

.PROBE TRAN
+    V(A)
+    V(B)
+    V(Cin)
+    V(S)

*.ALTER
** [0, 0] [0, 1]
*Vin1 A gnd 0v
*Vin2 B gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)

*.ALTER
** [0, 0] [1, 0]
*Vin1 A gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)
*Vin2 B gnd 0v

*.ALTER
** [0, 0] [1, 1]
*Vin1 A gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)
*Vin2 B gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)

*.ALTER
** [0, 1] [0, 0]
*Vin1 A gnd 0v
*Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)

*.ALTER
** [0, 1] [1, 1]  worst case!!
Vin1 A gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)
Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 9.8n 20n)
.MEASURE TRAN DELAY_COUT TRIG V(a) VAL=0.35 RISE=1 TARG V(COUT) VAL= 0.35 RISE=1
.MEASURE TRAN DELAY_S TRIG V(a) VAL=0.35 RISE=1 TARG V(S) VAL= 0.35 FALL=1

*.ALTER
** [1, 0] [0, 0]
*Vin1 A gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)
*Vin2 B gnd 0v

*.ALTER
** [1, 0] [1, 1]
*Vin1 A gnd PULSE (0v 0.7v 0n 0.1n 0.1n 9.8n 20n)
*Vin2 B gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 20n)

*.ALTER
** [1, 1] [0, 0]
*Vin1 A gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)
*Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)

*.ALTER
** [1, 1] [0, 1]
*Vin1 A gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)
*Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 9.8n 20n)

*.ALTER
** [1, 1] [1, 0]
*Vin1 A gnd PULSE (0v 0.7v 0n 0.1n 0.1n 9.8n 20n)
*Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 20n)


.END








