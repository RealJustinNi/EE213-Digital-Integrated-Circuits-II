*full adder
.TEMP 25
.OPTIONS ACCURATE
.OPTIONS POST=2

* YOU SHOULD INCLUDE MODLE FILES
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/NMOS_VTL.inc"
*.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/PMOS_VTL.inc"

* YOU SHOULD INCLUDE YOUR NELIST
.INCLUDE fulladder.sp

* YOU SHOULD ADD LOAD CAPACITANCE

* YOU SHOULD GIVE INPUT PATTERNS FOR TEST CASES
*Vin1 A gnd PULSE (0v 0.7v 19.9n 0.1n 0.1n 19.9n 40n)
*Vin2 B gnd PULSE (0v 0.7v 9.9n 0.1n 0.1n 9.9n 20n)
*Vin3 Cin gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 10n)

* YOU SHOULD GIVE PROPER INPUT PATTERNS FOR MAXIMUM DELAY

.PARAM PERIOD =40NS
.PARAM T0= 0.1NS
.PARAM T1= T0+PERIOD
.PARAM T2= T1+0.1NS
.PARAM STEP= 1PS

VDD   VDD! 0 0.7
VGND  GND! 0 0

.TRAN STEP T2

* YOU SHOULD MAKE SURE THAT YOU ARE MEASURING THE CORRECT SIGNAL FOR MAXIMUM DELAY. BELOW IS JUST AN EXAMPLE.
**[0 1 1]->[1 0 0 ]
Vin1 A gnd PULSE (0v 0.7v 4.9n 0.1n 0.1n 4.9n 40n)
Vin2 B gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 40n)
Vin3 Cin gnd PULSE (0v 0.7v 0n 0.1n 0.1n 4.9n 40n)
.MEASURE TRAN DELAY_COUT TRIG V(b) VAL=0.35 FALL=1 TARG V(COUT) VAL= 0.35 FALL=1
.MEASURE TRAN DELAY_S TRIG V(b) VAL=0.35 FALL=1 TARG V(S) VAL= 0.35 RISE=1

.PROBE TRAN
+    V(A)
+    V(B)
+    V(Cin)
+    V(Cout)
+    V(s)

.END








