** Generated for: hspiceD
** Generated on: Nov 13 20:51:14 2022
** Design library name: mylib2
** Design cell name: myHATestbench
** Design view name: schematic

.GLOBAL vdd!
.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/NMOS_VTL.inc"
.INCLUDE "/home/centos/PDK/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_ss/PMOS_VTL.inc"
.include "halfadder.pex.netlist.pex"

.subckt halfadder  A COUT S B GND! VDD!
* 
* VDD!	VDD!
* GND!	GND!
* B	B
* S	S
* COUT	COUT
* A	A
MM22 N_NET09_MM22_d N_A_MM22_g N_GND!_MM22_s N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=9e-08 AD=1.17e-14 AS=1.35e-14 PD=4.4e-07 PS=4.8e-07
MM25 N_NET07_MM25_d N_NET09_MM25_g N_GND!_MM22_s N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=9e-08 AD=1.08e-14 AS=1.35e-14 PD=4.2e-07 PS=4.8e-07
MM20 N_COUT_MM20_d N_NET14_MM20_g N_GND!_MM20_s N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=9e-08 AD=1.17e-14 AS=1.35e-14 PD=4.4e-07 PS=4.8e-07
MM0 N_NET14_MM0_d N_NET07_MM0_g NET056 N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM1 NET056 N_NET013_MM1_g N_GND!_MM1_s N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.7e-14 AS=2.16e-14 PD=6.6e-07 PS=6e-07
MM3 NET20 N_NET07_MM3_g N_GND!_MM3_s N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.7e-14 AS=2.34e-14 PD=6.6e-07 PS=6.2e-07
MM2 N_NET22_MM2_d N_NET14_MM2_g NET20 N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM19 N_S_MM19_d N_NET22_MM19_g NET35 N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM16 NET35 N_NET30_MM16_g N_GND!_MM16_s N_GND!_MM22_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.7e-14 AS=2.16e-14 PD=6.6e-07 PS=6e-07
MM12 N_NET30_MM12_d N_NET013_MM12_g NET055 N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM15 NET055 N_NET14_MM15_g N_GND!_MM15_s N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.7e-14 AS=2.16e-14 PD=6.6e-07 PS=6e-07
MM29 N_NET013_MM29_d N_NET017_MM29_g N_GND!_MM29_s N_GND!_MM22_b NMOS_VTL
+ L=5e-08 W=9e-08 AD=1.17e-14 AS=1.44e-14 PD=4.4e-07 PS=5e-07
MM26 N_NET017_MM26_d N_B_MM26_g N_GND!_MM29_s N_GND!_MM22_b NMOS_VTL L=5e-08
+ W=9e-08 AD=9.9e-15 AS=1.44e-14 PD=4e-07 PS=5e-07
MM23 N_NET09_MM23_d N_A_MM23_g N_VDD!_MM23_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM24 N_NET07_MM24_d N_NET09_MM24_g N_VDD!_MM23_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM21 N_COUT_MM21_d N_NET14_MM21_g N_VDD!_MM21_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM8 N_NET14_MM8_d N_NET07_MM8_g N_VDD!_MM8_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM9 N_NET14_MM9_d N_NET013_MM9_g N_VDD!_MM8_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM10 N_NET22_MM10_d N_NET07_MM10_g N_VDD!_MM10_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM11 N_NET22_MM11_d N_NET14_MM11_g N_VDD!_MM10_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM18 N_S_MM18_d N_NET22_MM18_g N_VDD!_MM18_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM17 N_S_MM17_d N_NET30_MM17_g N_VDD!_MM18_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM13 N_NET30_MM13_d N_NET013_MM13_g N_VDD!_MM13_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.34e-14 AS=2.7e-14 PD=6.2e-07 PS=6.6e-07
MM14 N_NET30_MM14_d N_NET14_MM14_g N_VDD!_MM13_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=2.16e-14 AS=2.7e-14 PD=6e-07 PS=6.6e-07
MM28 N_NET013_MM28_d N_NET017_MM28_g N_VDD!_MM28_s N_VDD!_MM23_b PMOS_VTL
+ L=5e-08 W=1.8e-07 AD=2.34e-14 AS=2.88e-14 PD=6.2e-07 PS=6.8e-07
MM27 N_NET017_MM27_d N_B_MM27_g N_VDD!_MM28_s N_VDD!_MM23_b PMOS_VTL L=5e-08
+ W=1.8e-07 AD=1.98e-14 AS=2.88e-14 PD=5.8e-07 PS=6.8e-07
*
.include "halfadder.pex.netlist.HALFADDER.pxi"
*
.ends
*
*

** Library name: mylib2
** Cell name: halfaddertb
** View name: schematic
xhalfadder a cout s b gnd! vdd! halfadder
c1 s 0 100e-15
c0 cout 0 100e-15


